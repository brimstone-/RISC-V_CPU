module sat_counter (
    input logic clk, 
    input logic [1:0] counter_val, 
    input logic do_count,       
    input logic is_count_up, 
    output logic [1:0] new_counter_val
);

endmodule: sat_counter 