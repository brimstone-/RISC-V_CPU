import rv32i_types::*;

module execute #(parameter width = 32)
(
	input clk,
	input stage_regs regs_in,
	output stage_regs regs_out
);

rv32i_word alumux1_out, alumux2_out;
rv32i_word cmpmux_out;

stage_regs regs;

logic br_en;

// ALU
mux2 alumux1
(
	.sel(regs_in.ctrl.alumux1_sel),
	.a(regs_in.rs1),
	.b(regs_in.pc),
	.f(alumux1_out)
);

mux8 alumux2
(
	.sel(regs_in.ctrl.alumux2_sel),
	.a(regs_in.i_imm),
	.b(regs_in.u_imm),
	.c(regs_in.b_imm),
	.d(regs_in.s_imm),
	.e(regs_in.rs2),
	.f(regs_in.j_imm),
	.g(),
	.h(),
	.out(alumux2_out)
);

alu alu
(
	.aluop(regs_in.ctrl.aluop),
	.a(alumux1_out),
	.b(alumux2_out),
	.f(regs_out.alu)
);

// CMP
mux2 cmpmux
(
	.sel(regs_in.ctrl.cmpmux_sel),
	.a(regs_in.rs2),
	.b(regs_in.i_imm),
	.f(cmpmux_out)
);

cmp cmp_module
(
	.cmpop(regs_in.ctrl.cmpop),
	.a(regs_in.rs1),
	.b(cmpmux_out),
	.br_en(br_en)
);

// stage_regs value passing
assign regs.i_imm = in.i_imm;
assign regs.s_imm = in.s_imm;
assign regs.b_imm = in.b_imm;
assign regs.u_imm = in.u_imm;
assign regs.j_imm = in.j_imm;
assign regs.rd = in.rd;
assign regs.rs1 = in.rs1;
assign regs.rs2 = in.rs2;
assign regs.pc = regs_out.alu;
assign regs.ctrl = in.ctrl;
assign regs.br = {{31{1'b0}},br_en};
assign regs.valid = in.valid;
assign regs.funct3 = in.funct3;

register #($bits(out)) stage_reg
(
	 .clk(clk),
    .load(1'b1), 					// always high for now. will be dependedent on mem_resp later
    .in(regs),						// struct of things to pass to stage 4
    .out(regs_out)						// values stage 3 holds
);

endmodule : execute
